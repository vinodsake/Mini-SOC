package my_pkg;
	parameter FIFO_DEPTH = 8;
	parameter DATA_WIDTH = 8;
endpackage
